
module PC_4 ( PC,PCN);
input [31:0] PC;
output [31:0] PCN ;

assign PCN=PC + 4;


		
endmodule 
